module m1;

global int exportedVar = 42;
global int otherVar = 4242;
