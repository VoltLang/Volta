//T compiles:yes
//T retval:12
// Combining addition and subtraction.
module test_003;

int main()
{
    return 12 - 6 + 12 - 6;
}
