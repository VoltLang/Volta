//T compiles:no
module test_017;

int main()
{
	string foo = 4;

	return 42;
}
