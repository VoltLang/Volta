module m8;

import ctx = m1;
