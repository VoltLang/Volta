//T compiles:yes
//T retval:78
// Simple subtraction.
module test_002;

int main()
{
    return 82 - 4;
}
