//T compiles:no
// Test appending to an array, expected to fail.

module test_018;

int main()
{
	short[] s;
	int i = 3;
	s ~= i;
}
