//T compiles:yes
//T retval:32
// Local var test.
module test_003;

local int var;

int main()
{
	var = 32;
	return var;
}
