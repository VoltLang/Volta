//T compiles:yes
//T retval:16
// Parens and order of evaluation.
module test_005;

int main()
{
    return 4 * (5 - 1);
}
