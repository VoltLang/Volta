//T compiles:yes
//T retval:42
// Most basic test.
module test_001;

int main()
{
	return 42;
}
