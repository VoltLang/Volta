//T compiles:yes
//T retval:16
// Hexadecimal literals.
module test_011;

int main()
{
    return 0x10;
}
