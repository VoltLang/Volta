//T compiles:yes
//T retval:1
// Condition to bool.
module test_017;

int main()
{
	return 1 ? 1 : 2;
}
